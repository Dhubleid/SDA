library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package Matrix is    

type mat is array(natural range <>) of std_logic_vector(7 downto 0);
	
end Matrix;

